// Build a circuit with no inputs and one output that outputs a constant 0
module top_module (
    output zero
    // not assigning a value to a signal usually results in 0
);
  
endmodule
