// learn the use with assign
// "assign a = b" mean copy b value to a
module top_module( input in, output out );
    assign out = in;
endmodule
