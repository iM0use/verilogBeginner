module top_module( output one );
    // Build a circuit with no inputs and one output. That output should always drive 1 (or logic high). 
    assign one = 1;
endmodule
